module cxf
