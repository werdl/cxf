module main

import cxf

fn main() {
	fifty := cxf.cxf('-50')
	println(cxf.pad('76835874', 6))
}
