module main

import cxf

fn main() {
	fifty := cxf.cxf('50')
	println(fifty.bin())
}
